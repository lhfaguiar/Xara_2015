-- Arquivo maior (?)
-- 20151209
--

-- ------------------------------------
--  THE XARA PROJECT
-- ------------------------------------
--  Author : Lai Aguiar
---------------------------------------



library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity Xara_20151209 is
    port(

    );
end Xara_20151209;

-- architecture Xara of Xara_20151209 is

--     component Xara_DF
--         port(
--             progr                           : in std_logic_vector (15 downto 0);
--             memoria                         : out std_logic_vector (15 downto 0);
--             S                               : in std_logic_vector(3 downto 0);
--             CIN, R1, R0                     : in std_logic_vector (1 downto 0);
--             grava, clear_4regs              : in std_logic;
--             decoder_en, neg_clear_counter   : in std_logic;
--             count_en, load_reg_saida        : in std_logic;
--             R20, R21                        : in std_logic;
--             CLOCK                           : in std_logic;
--             CLEAR                           : in std_logic;
--             modo_memoria                    : in std_logic;
--             modo_mem                        : out std_logic;
--             limpa                           : in std_logic;
--             limpa_s                         : out std_logic
--         );
--     end component;

--     component Xara_cu
--         port(

--         );
--     end component;


    -- sinais!!

    -- controlunit
    -- Xara_cu : controlunit
    --     portmap (
    --         memoria             =>
    --         S                   =>
    --         CIN                 =>
    --         R1                  =>
    --         R0                  =>
    --         grava               =>
    --         clear_4regs         =>
    --         decoder_en          =>
    --         neg_clear_counter   =>
    --         count_en            =>
    --         load_reg_saida      =>
    --         R20, R21            =>
    --         CLOCK               =>
    --         CLEAR               =>
    --         modo_memoria        =>
    --     );

    -- Xara_DF : data_flow
    --     portmap (

    --     );
